module Hello;
initial
begin : main

	$display ("Hello World!");

end
endmodule
	
